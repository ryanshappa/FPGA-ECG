library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
  
entity ShiftR is
port ( 
	
end ADCClk;
  
architecture behavior of ShiftR is